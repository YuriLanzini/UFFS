module registrador();

endmodule
